module Hazard_Detection(
    Stall_o
);

output Stall_o;

assign Stall_o = 0;

endmodule